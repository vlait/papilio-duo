-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity DECODER_6 is
port (
	CLK  : in  std_logic;
	ADDR : in  std_logic_vector(8 downto 0);
	DATA : out std_logic_vector(7 downto 0);
	DI   : in std_logic_vector(7 downto 0);
	WE   : in std_logic
	);
end;

architecture RTL of DECODER_6 is

	signal rom_addr : std_logic_vector(10 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(8 downto 0) <= ADDR;
	end process;

	DECODER_6_0 : RAMB16_S9
	generic map (
		INITP_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => x"0000000000000000000000000000000000000000000000000000000000000000",

		INIT_00 => x"1E1D1C1B1A191817161514131211100F0E0D0C0B0A0908070605040302010000",
		INIT_01 => x"3E3D3C3B3A393837363534333231302F2E2D2C2B2A292827262524232221201F",
		INIT_02 => x"5E5D5C5B5A595857565554535251504F4E4D4C4B4A494847464544434241403F",
		INIT_03 => x"7E7D7C7B7A797877767574737271706F6E6D6C6B6A696867666564636261605F",
		INIT_04 => x"9E9D9C9B9A999897969594939291908F8E8D8C8B8A898887868584838281807F",
		INIT_05 => x"BEBDBCBBBAB9B8B7B6B5B4B3B2B1B0AFAEADACABAAA9A8A7A6A5A4A3A2A1A09F",
		INIT_06 => x"DEDDDCDBDAD9D8D7D6D5D4D3D2D1D0CFCECDCCCBCAC9C8C7C6C5C4C3C2C1C0BF",
		INIT_07 => x"00000000000000F7F6F5F4F3F2F1F0EFEEEDECEBEAE9E8E7E6E5E4E3E2E1E0DF",
		INIT_08 => x"DFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F700000000000000",
		INIT_09 => x"BFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDE",
		INIT_0A => x"9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBE",
		INIT_0B => x"7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E",
		INIT_0C => x"5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E",
		INIT_0D => x"3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E",
		INIT_0E => x"1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E",
		INIT_0F => x"00000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 0),
		DOP  => open,
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => DI,
--		DI   => "00000000",
		DIP  => "0",
		EN   => '1',
		SSR  => '0',
		WE   => WE
--		WE   => '0'
	);

end RTL;
