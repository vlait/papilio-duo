-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity DECODER_4 is
port (
	CLK  : in  std_logic;
	ADDR : in  std_logic_vector(8 downto 0);
	DATA : out std_logic_vector(7 downto 0);
	DI   : in std_logic_vector(7 downto 0);
	WE   : in std_logic
	);
end;

architecture RTL of DECODER_4 is

	signal rom_addr : std_logic_vector(10 downto 0);

begin

	p_addr : process(ADDR)
	begin
		rom_addr <= (others => '0');
		rom_addr(8 downto 0) <= ADDR;
	end process;

	DECODER_4_0 : RAMB16_S9
	generic map (
		INITP_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => x"0000000000000000000000000000000000000000000000000000000000000000",

		INIT_00 => x"0C8B4B0B8A4A0A89490988480887470786460685450584440483430382420281",
		INIT_01 => x"9656169555159454149353139252129151119050108F4F0F8E4E0E8D4D0D8C4C",
		INIT_02 => x"6121A060209F5F1F9E5E1E9D5D1D9C5C1C9B5B1B9A5A1A995919985818975717",
		INIT_03 => x"2CAB6B2BAA6A2AA96929A86828A76727A66626A56525A46424A36323A26222A1",
		INIT_04 => x"B67636B57535B47434B37333B27232B17131B07030AF6F2FAE6E2EAD6D2DAC6C",
		INIT_05 => x"4101804000BF7F3FBE7E3EBD7D3DBC7C3CBB7B3BBA7A3AB97939B87838B77737",
		INIT_06 => x"C3C5CCC580D3CDC1C9CCCCC9D780B1B8B9B180A9C3A880D4C8C7C9D2D9D0CFC3",
		INIT_07 => x"C4C5D6D2C5D3C5D280D3D4C8C7C9D280CCCCC180AEC3CEC980D3C3C9CECFD2D4",
		INIT_08 => x"A92A6AAA2B6BAB2C6CAC2D6DAD2E6EAE2F6FAF3070B03171B13272B23373B334",
		INIT_09 => x"1F5F9F2060A02161A12262A22363A32464A42565A52666A62767A72868A82969",
		INIT_0A => x"54941555951656961757971858981959991A5A9A1B5B9B1C5C9C1D5D9D1E5E9E",
		INIT_0B => x"890A4A8A0B4B8B0C4C8C0D4D8D0E4E8E0F4F8F10509011519112529213539314",
		INIT_0C => x"B67636B57535B474810242820343830444840545850646860747870848880949",
		INIT_0D => x"4101804000BF7F3FBE7E3EBD7D3DBC7C3CBB7B3BBA7A3AB97939B87838B77737",
		INIT_0E => x"C3C5CCC580D3CDC1C9CCCCC9D780B1B8B9B180A9C3A880D4C8C7C9D2D9D0CFC3",
		INIT_0F => x"C4C5D6D2C5D3C5D280D3D4C8C7C9D280CCCCC180AEC3CEC980D3C3C9CECFD2D4",
		INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DO   => DATA(7 downto 0),
		DOP  => open,
		ADDR => rom_addr,
		CLK  => CLK,
		DI   => DI,
--		DI   => "00000000",
		DIP  => "0",
		EN   => '1',
		SSR  => '0',
		WE	  => WE
--		WE   => '0'
	);

end RTL;
